module processing_block (
  left_input, middle_input, right_input,
  left_output, middle_output, right_output,
  filter_output
)
  // Reg: have 3x3 reg, that on ready shifts all data upward by one



endmodule
